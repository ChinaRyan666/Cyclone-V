module  FullConnect_WriteBuffer #(
    parameter                       AvalonData_WIDTH        =   512
)  (

    //  General Signals
    input   wire                clk,
    input   wire                rstn,

    //  From Piplined MAC
    input   wire                Valid_i,
    output  wire                Halt_o,
    input   wire    [31:0]      Data_i,
    
    //  To WriteMaster
    output  wire    [AvalonData_WIDTH-1:0]     WriteData_o,
    output  wire                WriteReq_o,
    input   wire                WriteAck_i

);



//  WRITEBUFFER TAG
wire      BufferWrite;
wire[31:0]      Data_ireg;

assign  BufferWrite  = Valid_i &   ~Halt_o;


FullConnectDFF #(
    .WIDTH      (1),
    .RstVal     (1'b0),
    .PstVal     (1'b0)
)   WriteBufferTag (
    .clk        (clk),
    .rstn       (rstn),
    .Set_i      (WriteAck_i & WriteReq_o),
    .Enable_i   (BufferWrite),
    .D_i        (1'b1),
    .Q_o        (WriteReq_o)
);

FullConnectDFF #(
    .WIDTH      (32),
    .RstVal     (1'b0),
    .PstVal     (1'b0)
)   DataTag (
    .clk        (clk),
    .rstn       (rstn),
    .Set_i      (1'b0),
    .Enable_i   (1'b1),
    .D_i        (Data_i),
    .Q_o        (Data_ireg)
);
assign WriteData_o = {{(AvalonData_WIDTH-32){1'b0}},Data_ireg};

assign  Halt_o  =   WriteReq_o & Valid_i;



endmodule